LIBRARY ieee;
USE IEEE.std_logic_1164.ALL;

LIBRARY work;

PACKAGE ASCII IS
  SUBTYPE ASCII IS std_logic_vector(7 DOWNTO 0);

  CONSTANT A : ASCII := "01000001";
  CONSTANT B : ASCII := "01000010";
  CONSTANT C : ASCII := "01000011";
  CONSTANT D : ASCII := "01000100";
  CONSTANT E : ASCII := "01000101";
  CONSTANT F : ASCII := "01000110";
  CONSTANT G : ASCII := "01000111";
  CONSTANT H : ASCII := "01001000";
  CONSTANT I : ASCII := "01001001";
  CONSTANT J : ASCII := "01001010";
  CONSTANT K : ASCII := "01001011";
  CONSTANT L : ASCII := "01001100";
  CONSTANT M : ASCII := "01001101";
  CONSTANT N : ASCII := "01001110";
  CONSTANT O : ASCII := "01001111";
  CONSTANT P : ASCII := "01010000";
  CONSTANT Q : ASCII := "01010001";
  CONSTANT R : ASCII := "01010010";
  CONSTANT S : ASCII := "01010011";
  CONSTANT T : ASCII := "01010100";
  CONSTANT U : ASCII := "01010101";
  CONSTANT V : ASCII := "01010110";
  CONSTANT W : ASCII := "01010111";
  CONSTANT X : ASCII := "01011000";
  CONSTANT Y : ASCII := "01011001";
  CONSTANT Z : ASCII := "01011010";

  CONSTANT d0 : ASCII := "00110000";
  CONSTANT d1 : ASCII := "00110001";
  CONSTANT d2 : ASCII := "00110010";
  CONSTANT d3 : ASCII := "00110011";
  CONSTANT d4 : ASCII := "00110100";
  CONSTANT d5 : ASCII := "00110101";
  CONSTANT d6 : ASCII := "00110110";
  CONSTANT d7 : ASCII := "00110111";
  CONSTANT d8 : ASCII := "00111000";
  CONSTANT d9 : ASCII := "00111001";
END;