LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY CallPlatform IS
  PORT (
    clock : IN std_logic
    -- TODO
  );
END CallPlatform;

ARCHITECTURE rtl OF CallPlatform IS
  -- TODO
BEGIN
  -- TODO
END rtl;