LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.ALL;

LIBRARY work;
USE work.config.ALL;

-- ����Դ -> ȡ�� -> ���� -> ������
ENTITY Service IS
  PORT (
    clock : IN std_logic;
    reset : IN std_logic;
    call : IN std_logic; -- �к�
    recall : IN std_logic; -- ���½к�

    pull : OUT std_logic; -- ����ȡ��
    empty : IN std_logic; -- ����Ϊ��
    enable_pull : IN std_logic; -- ����ȡ��

    push : OUT std_logic; -- ���뷢��
    pushed : IN std_logic; -- �ѷ���

    data_in : IN std_logic_vector(RAM_WIDTH - 1 DOWNTO 0);
    data_out : OUT std_logic_vector(RAM_WIDTH - 1 DOWNTO 0)
  );
END Service;

ARCHITECTURE arch OF Service IS
  TYPE states IS(idle, start, queue_empty, pulling, pushing);
  SIGNAL present_state : states;
  SIGNAL next_state : states;

  SIGNAL data : std_logic_vector(RAM_WIDTH - 1 DOWNTO 0);
  CONSTANT DATA_DEFAULT : std_logic_vector(DATA_WIDTH - 1 DOWNTO 0) := (OTHERS => '0');

  -- jump next state
  FUNCTION ifElse(
    condition : std_logic;
    onTrue : states;
    onFalse : states
  ) RETURN states IS
  BEGIN
    IF (condition = '1') THEN
      RETURN onTrue;
    ELSE
      RETURN onFalse;
    END IF;
  END FUNCTION;
BEGIN
  -- clock trigger
  PROCESS (clock, reset)
  BEGIN
    IF (reset = '1') THEN
      present_state <= idle;
    ELSIF (clock'event AND clock = '1') THEN
      present_state <= next_state;
    END IF;
  END PROCESS;

  -- state change
  PROCESS (present_state, call, recall, enable_pull, empty, pushed)
  BEGIN
    CASE present_state IS
      WHEN idle =>
        IF (call = '1') THEN
          next_state <= pulling;
        ELSIF (recall = '1') THEN
          next_state <= pushing;
        ELSE
          next_state <= idle;
        END IF;

      WHEN start =>
        next_state <= ifElse(empty, queue_empty, pulling);

      WHEN queue_empty =>
        next_state <= pushing;

      WHEN pulling =>
        next_state <= ifElse(enable_pull, pushing, pulling);

      WHEN pushing =>
        next_state <= ifElse(pushed, idle, pushing);

      WHEN OTHERS =>
        next_state <= idle;
    END CASE;
  END PROCESS;

  -- state events
  PROCESS (present_state, data_in, data)
  BEGIN
    -- make latches: data
    push <= '0';
    pull <= '0';
    data_out <=
      FLAG_SCREEN_SERVICE &
      FLAG_ERROR_UNKNOWN &
      FLAG_GROUP_FREE &
      DATA_DEFAULT;

    CASE present_state IS
      WHEN idle => NULL;

      WHEN pulling =>
        pull <= '1';
        data <=
          FLAG_SCREEN_SERVICE &
          data_in(FLAG_SCREEN_LOW - 1 DOWNTO 0);

      WHEN queue_empty =>
        data <=
          FLAG_SCREEN_SERVICE &
          FLAG_ERROR_QUEUE_EMPTY &
          data(FLAG_GROUP_HIGH DOWNTO 0);

      WHEN pushing =>
        push <= '1';
        data_out <= data;

      WHEN OTHERS => NULL;

    END CASE;
  END PROCESS;
END arch;